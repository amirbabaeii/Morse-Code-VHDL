---- fpga4student.com: FPGA projects, Verilog projects, VHDL projects 
---- VHDL project: VHDL code for a single-port RAM 
--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;
--USE ieee.numeric_std.ALL;
--
---- A 128x8 single-port RAM in VHDL
--entity Single_port_RAM_VHDL is
--port(
-- RAM_ADDR: in integer range 0 to 607; -- Address to write/read RAM
-- RAM_DATA_IN: in std_logic_vector(0 to 7); -- Data to write into RAM
-- RAM_WR: in std_logic; -- Write enable 
-- RAM_CLOCK: in std_logic; -- clock input for RAM
-- RAM_DATA_OUT: out std_logic_vector(0 to 7) -- Data output of RAM
--);
--end Single_port_RAM_VHDL;
--
--architecture Behavioral of Single_port_RAM_VHDL is
---- define the new type for the 128x8 RAM 
--type RAM_ARRAY is array (0 to 607,0 to 7) of std_logic;
---- initial values in the RAM
--signal RAM: RAM_ARRAY :=(
--				"00000000",
--				"00000000",
--				"00010000",
--				"00111000",
--				"01101100",
--				"11000110",
--				"11000110",
--				"11111110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- A ---
--				"00000000",
--				"00000000",
--				"11111000",
--				"11001100",
--				"11000110",
--				"11001100",
--				"11111100",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11001100",
--				"11111000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- B ---
--				"00000000",
--				"00000000",
--				"01111100",
--				"11001110",
--				"11000110",
--				"11000000",
--				"11000000",
--				"11000000",
--				"11000000",
--				"11000110",
--				"11001110",
--				"01111100",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- C ---
--				"00000000",
--				"00000000",
--				"11111000",
--				"11001100",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11001100",
--				"11111000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- D ---
--				"00000000",
--				"00000000",
--				"11111110",
--				"11000010",
--				"11000000",
--				"11000100",
--				"11111100",
--				"11000100",
--				"11000000",
--				"11000000",
--				"11000010",
--				"11111110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- E ---
--				"00000000",
--				"00000000",
--				"11111110",
--				"11000010",
--				"11000000",
--				"11000100",
--				"11111100",
--				"11000100",
--				"11000000",
--				"11000000",
--				"11000000",
--				"11100000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- F ---
--				"00000000",
--				"00000000",
--				"11111110",
--				"11000110",
--				"11000010",
--				"11000000",
--				"11000000",
--				"11001110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11111110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- G ---
--				"00000000",
--				"00000000",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11111110",
--				"11111110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- H ---
--				"00000000",
--				"00000000",
--				"00111100",
--				"00011000",
--				"00011000",
--				"00011000",
--				"00011000",
--				"00011000",
--				"00011000",
--				"00011000",
--				"00011000",
--				"00111100",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- I ---
--				"00000000",
--				"00000000",
--				"00011110",
--				"00001100",
--				"00001100",
--				"00001100",
--				"00001100",
--				"00001100",
--				"00001100",
--				"11001100",
--				"11001100",
--				"01111000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- J ---
--				"00000000",
--				"00000000",
--				"11000110",
--				"11001100",
--				"11011000",
--				"11110000",
--				"11100000",
--				"11110000",
--				"11011000",
--				"11001100",
--				"11000110",
--				"11000010",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- K ---
--				"00000000",
--				"00000000",
--				"11000000",
--				"11000000",
--				"11000000",
--				"11000000",
--				"11000000",
--				"11000000",
--				"11000000",
--				"11000000",
--				"11000110",
--				"11111110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- L ---
--				"00000000",
--				"00000000",
--				"11101110",
--				"10101010",
--				"10101010",
--				"10101010",
--				"10111010",
--				"10010010",
--				"10000010",
--				"10000010",
--				"10000010",
--				"10000010",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- M ---
--				"00000000",
--				"00000000",
--				"11100010",
--				"10100010",
--				"10100010",
--				"10100010",
--				"10010010",
--				"10010010",
--				"10010010",
--				"10001010",
--				"10001010",
--				"10001110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- N ---
--				"00000000",
--				"00000000",
--				"00111000",
--				"01101100",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"01101100",
--				"00111000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- O ---
--				"00000000",
--				"00000000",
--				"11111000",
--				"11001100",
--				"11000110",
--				"11000110",
--				"11001110",
--				"11111000",
--				"11000000",
--				"11000000",
--				"11000000",
--				"11100000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- P ---
--				"00000000",
--				"00000000",
--				"00111000",
--				"01101100",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11010110",
--				"01101100",
--				"00111010",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- Q ---
--				"00000000",
--				"00000000",
--				"11111000",
--				"11001100",
--				"11000110",
--				"11000110",
--				"11001110",
--				"11111000",
--				"11110000",
--				"11011000",
--				"11001100",
--				"11000110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- R ---
--				"00000000",
--				"00000000",
--				"01111110",
--				"11000000",
--				"11000000",
--				"01100000",
--				"00110000",
--				"00011000",
--				"00001100",
--				"00000110",
--				"00001100",
--				"11111000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- S ---
--				"00000000",
--				"00000000",
--				"11111110",
--				"10010010",
--				"00010000",
--				"00010000",
--				"00010000",
--				"00010000",
--				"00010000",
--				"00010000",
--				"00010000",
--				"00111000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- T ---
--				"00000000",
--				"00000000",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"01101100",
--				"00111000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- U ---
--				"00000000",
--				"00000000",
--				"11000110",
--				"11000110",
--				"11000110",
--				"01101100",
--				"01101100",
--				"01101100",
--				"00111000",
--				"00111000",
--				"00010000",
--				"00010000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- V ---
--				"00000000",
--				"00000000",
--				"10000010",
--				"10000010",
--				"10000010",
--				"10000010",
--				"10111010",
--				"10101010",
--				"10101010",
--				"10101010",
--				"10101010",
--				"11101110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- W ---
--				"00000000",
--				"00000000",
--				"11000110",
--				"11000110",
--				"01101100",
--				"01101100",
--				"00111000",
--				"01111100",
--				"01101100",
--				"01101100",
--				"11000110",
--				"11000110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- X ---
--				"00000000",
--				"00000000",
--				"11000110",
--				"11000110",
--				"11000110",
--				"01101100",
--				"00111000",
--				"00010000",
--				"00010000",
--				"00010000",
--				"00010000",
--				"00010000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- Y ---
--				"00000000",
--				"00000000",
--				"11111110",
--				"11111110",
--				"00000110",
--				"00001100",
--				"00011000",
--				"00110000",
--				"01100000",
--				"11000000",
--				"11111110",
--				"11111110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- Z ---
--				"00000000",
--				"00000000",
--				"01111100",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"01111100",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- ZERO ---
--				"00000000",
--				"00000000",
--				"00111000",
--				"01011000",
--				"00011000",
--				"00011000",
--				"00011000",
--				"00011000",
--				"00011000",
--				"00011000",
--				"00111100",
--				"00111100",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- ONE ---
--				"00000000",
--				"00000000",
--				"11111100",
--				"11000110",
--				"11000110",
--				"00001100",
--				"00011000",
--				"00110000",
--				"11000000",
--				"11000000",
--				"11111110",
--				"11111110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- TWO ---
--				"00000000",
--				"00000000",
--				"01111100",
--				"11000110",
--				"01000110",
--				"00000110",
--				"00000100",
--				"00111100",
--				"00000100",
--				"01000110",
--				"11000110",
--				"01111100",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- THREE ---
--				"00000000",
--				"00000000",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11000110",
--				"11111110",
--				"11111110",
--				"00000110",
--				"00000110",
--				"00000110",
--				"00000110",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- FOUR ---
--				"00000000",
--				"00000000",
--				"11111110",
--				"11111110",
--				"11000000",
--				"11000000",
--				"01110000",
--				"00011000",
--				"00001100",
--				"00000110",
--				"11001100",
--				"11111000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- FIVE ---
--				"00000000",
--				"00000000",
--				"00000110",
--				"00001100",
--				"00011000",
--				"00110000",
--				"01100000",
--				"11111100",
--				"11000110",
--				"11000110",
--				"01100110",
--				"00111100",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- SIX ---
--				"00000000",
--				"00000000",
--				"11111110",
--				"11111100",
--				"00001100",
--				"00011000",
--				"00011000",
--				"00110000",
--				"00110000",
--				"01100000",
--				"01100000",
--				"11000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- SEVEN ---
--				"00000000",
--				"00000000",
--				"00111000",
--				"01101100",
--				"11000110",
--				"01101100",
--				"00111000",
--				"01101100",
--				"11000110",
--				"11000110",
--				"01101100",
--				"00111000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- EIGHT ---
--				"00000000",
--				"00000000",
--				"00111100",
--				"01100110",
--				"11000110",
--				"11000110",
--				"01100110",
--				"00111110",
--				"00000110",
--				"00000110",
--				"00001100",
--				"11111000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- NINE ---
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000", --- SPACE ---
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00011000",
--				"00011000",
--				"00000000",
--				"00000000",
--				"00000000",
--				"00000000" --- DOT ---
--);
--begin
--process(RAM_CLOCK)
--begin
-- if(rising_edge(RAM_CLOCK)) then
-- if(RAM_WR='1') then -- when write enable = 1, 
-- -- write input data into RAM at the provided address
-- RAM(RAM_ADDR) <= RAM_DATA_IN;
-- -- The index of the RAM array type needs to be integer so
-- -- converts RAM_ADDR from std_logic_vector -> Unsigned -> Interger using numeric_std library
-- end if;
-- end if;
--end process;
-- -- Data to be read out 
-- RAM_DATA_OUT <= RAM(RAM_ADDR);
--end Behavioral;